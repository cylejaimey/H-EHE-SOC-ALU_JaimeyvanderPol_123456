--------------------------------------------------------------------
--! \file      sevenOut4Decoder.vhd
--! \date      11-1-2021
--! \brief     Place holder
--! \author    Remko Welling (WLGRW) remko.welling@han.nl
--! \copyright HAN TF ELT/ESE Arnhem 
------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.all;
------------------------------------------------------------------------------
ENTITY sevenOut4Decoder is

   PORT (
      input   : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
      dot     : IN  STD_LOGIC;
      ctrl    : IN  STD_LOGIC;
      display : OUT STD_LOGIC_VECTOR(0 TO 7)
   );
   
END ENTITY sevenOut4Decoder;
------------------------------------------------------------------------------
ARCHITECTURE implementation OF sevenOut4Decoder IS
BEGIN

--  #########################################################################
--  #########################################################################
--  ##                                                                     ##
--  ##                                                                     ##
--  ##  This file shall be replaced by the file produced in assignment 2-1 ##
--  ##                                                                     ##
--  ##                                                                     ##
--  #########################################################################
--  #########################################################################


END ARCHITECTURE implementation;
------------------------------------------------------------------------------
